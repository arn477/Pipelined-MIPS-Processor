library verilog;
use verilog.vl_types.all;
entity ALUControlUnit_vlg_vec_tst is
end ALUControlUnit_vlg_vec_tst;
