module CPU (clk, reset);
endmodule
