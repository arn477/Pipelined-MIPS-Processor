library verilog;
use verilog.vl_types.all;
entity signExtend_vlg_vec_tst is
end signExtend_vlg_vec_tst;
