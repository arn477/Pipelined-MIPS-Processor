//supports 15 instructions of 32 bit size
module InstructionMem(instruction, address);
	output [31:0] instruction;
	input [31:0] address;
	wire [3:0] rom_addr;
	reg[31:0] rom[14:0];

	
	assign rom_addr[3:0] = address[5:2];
	
	initial begin
		rom[0] = 32'b00111000000100000000000000000011;
		rom[1] = 32'b00111000000100010000000000000100;
		rom[2] = 32'b00001000000000000000000000000101;
		rom[3] = 32'b00111000000100000000000000000001;
		rom[4] = 32'b00111000000100010000000000000001;
		rom[5] = 32'b00000010001100001001000000100010;
		rom[6] = 32'b00010110000100011111111111111100;
		rom[7] = 32'b00000010000100011001100000100000;
		rom[8] = 32'b10101110010100110000000000010000;
		rom[9] = 32'b10001110010101000000000000010000;
		rom[10] = 32'b00000010000101001010100000101010;
		rom[11] = 32'b10001110010100110000000000010000;
		rom[12] = 32'b00111010010100110000000000000001;
		rom[13] = 32'b00111010101101010000000000000001;
		rom[14] = 32'b00000010101000000000000000001000;
	end
	
	assign instruction = (address[31:0]<60)?rom[rom_addr[3:0]]:32'd0;

endmodule
	