`timescale 1 ps / 100 fs
//supports 15 instructions of 32 bit size
module InstructionMem(instruction, address);
	output [31:0] instruction;
	input [31:0] address;
	wire [3:0] rom_addr;
	reg[31:0] rom[14:0];

	
	assign rom_addr[3:0] = address[5:2];
	
	initial begin
		rom[0] = 32'b00100000000100010000000000000001;
		rom[1] = 32'b00100000000100100000000000000010;
		rom[2] = 32'b00100000000100110000000000000011;
		rom[3] = 32'b00000010011100011010000000100000;
		rom[4] = 32'b00100010100101010000000000000010;
		rom[5] = 32'b00101010101010100000000000001010;
		rom[6] = 32'b10101110110101010000000000001000;
		rom[7] = 32'b00010010001010100000000000000001;
		rom[8] = 32'b00100010001100100000000000000100;
		rom[9] = 32'b00000010001100100100000000100101;
		rom[10] = 32'b00001000000000000000000000001100;
		rom[11] = 32'b00100000000010010000000000100000;
		rom[12] = 32'b10001110110100000000000000001000;
		rom[13] = 32'b00000000000000000000000000000000;
		rom[14] = 32'b00000000000000000000000000000000;
	end
	
	assign instruction = (address[31:0]<60)?rom[rom_addr[3:0]]:32'd0;

endmodule
	